
`include "global.v"


module bias_conv1_rom(
	input							clk,
	input							rst_n,
	input	[6:0]					aa,
	input							cena,
	output reg	[`WD_BIAS*4 -1:0]	qa
	);
	
	logic [0:0][0:3][`WD_BIAS-1:0] weight	 = {	
-12'd199,  12'd715,  -12'd124,  -12'd198
	};
	


	always @(posedge clk or negedge rst_n)
		if (!rst_n)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule

module wieght_conv1_rom(
	input						clk,
	input						rst_n,
	input	[9:0]				aa,
	input						cena,
	output reg	[`WD*4 -1:0]	qa
	);
	
	
	logic [0:24][0:3][`WD-1:0] weight	 = {
-8'd48,  -8'd83,  8'd43,  8'd75,  
-8'd56,  -8'd72,  8'd16,  8'd69,  
8'd35,  -8'd104,  -8'd5,  8'd22,  
8'd86,  -8'd85,  -8'd5,  -8'd41,  
8'd70,  -8'd71,  -8'd35,  -8'd80,  

-8'd117,  -8'd117,  8'd51,  8'd56,  
-8'd8,  -8'd85,  8'd7,  8'd91,  
8'd62,  -8'd60,  -8'd4,  8'd90,  
8'd74,  -8'd53,  -8'd19,  8'd20,  
8'd17,  -8'd90,  8'd21,  -8'd54,  

-8'd96,  -8'd81,  8'd68,  -8'd45,  
8'd63,  -8'd45,  8'd32,  8'd47,  
8'd85,  -8'd27,  8'd48,  8'd106,  
8'd94,  8'd20,  8'd38,  8'd76,  
-8'd67,  -8'd6,  8'd71,  -8'd13,  

-8'd13,  8'd57,  8'd79,  -8'd126,  
8'd60,  8'd90,  8'd47,  -8'd26,  
8'd85,  8'd101,  8'd42,  8'd59,  
8'd17,  8'd73,  8'd63,  8'd83,  
-8'd65,  8'd49,  8'd71,  8'd44,  

8'd61,  8'd109,  8'd32,  -8'd85,  
8'd63,  8'd63,  8'd39,  -8'd69,  
8'd30,  8'd50,  8'd31,  -8'd57,  
8'd5,  8'd23,  8'd6,  8'd48,  
-8'd34,  8'd61,  8'd26,  8'd59
		};

//5*5*4*8

	always @(posedge clk or negedge rst_n)
		if (!rst_n)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
	


endmodule	



module bias_fc1_rom(
	input							clk,
	input							rst_n,
	input	[6:0]					aa,
	input							cena,
	output reg	[`WD_BIAS*1 -1:0]	qa
	);
	
	logic [0:9][`WD_BIAS-1:0] weight	 = {
12'd167,  12'd485,  -12'd61,  -12'd432,  12'd111,  12'd219,  -12'd68,  12'd412,  -12'd518,  -12'd253	
	};
	
//120*1*24

	always @(posedge clk or negedge rst_n)
		if (!rst_n)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule

module wieght_fc1_rom(
	input							clk,
	input							rst_n,
	input	[11:0]					aa,
	input							cena,
	output reg	[`WD*4*1 -1:0]	qa
	);
	


	logic [0:10*7*7-1][0:3][`WD-1:0] weight	 = {
8'd8,  -8'd8,  -8'd18,  -8'd26,  8'd3,  8'd5,  -8'd3,  
-8'd1,  8'd0,  8'd12,  8'd6,  -8'd11,  8'd20,  -8'd17,  
-8'd15,  -8'd4,  -8'd14,  8'd9,  -8'd26,  8'd4,  -8'd10,  
-8'd8,  -8'd5,  -8'd4,  -8'd25,  8'd14,  8'd0,  -8'd28,  
-8'd11,  8'd11,  -8'd2,  -8'd13,  8'd7,  -8'd3,  8'd3,  
-8'd20,  -8'd13,  -8'd27,  -8'd27,  -8'd18,  -8'd1,  8'd8,  
8'd9,  8'd16,  -8'd8,  8'd6,  -8'd4,  8'd10,  8'd1,  
-8'd7,  8'd6,  -8'd7,  -8'd27,  -8'd4,  8'd28,  -8'd21,  
-8'd11,  8'd1,  -8'd24,  -8'd18,  8'd12,  8'd1,  8'd9,  
-8'd20,  8'd16,  -8'd1,  8'd6,  8'd22,  8'd18,  -8'd26,  
-8'd19,  8'd1,  -8'd29,  -8'd53,  -8'd6,  8'd59,  8'd4,  
-8'd54,  8'd27,  8'd22,  8'd15,  -8'd4,  8'd9,  -8'd30,  
-8'd32,  -8'd8,  -8'd7,  8'd4,  8'd25,  -8'd3,  8'd25,  
-8'd14,  8'd47,  -8'd33,  -8'd19,  -8'd10,  -8'd15,  -8'd56,  
-8'd54,  -8'd45,  8'd13,  -8'd31,  -8'd31,  -8'd5,  8'd32,  
-8'd41,  8'd15,  -8'd5,  8'd22,  -8'd59,  8'd39,  8'd35,  
-8'd14,  8'd14,  8'd19,  -8'd8,  8'd28,  -8'd81,  -8'd6,  
-8'd3,  8'd43,  -8'd59,  8'd21,  -8'd3,  -8'd21,  8'd27,  
8'd8,  -8'd15,  8'd15,  8'd4,  8'd17,  -8'd38,  8'd11,  
-8'd35,  8'd25,  8'd3,  8'd0,  -8'd41,  8'd34,  8'd18,  
8'd3,  -8'd25,  8'd19,  8'd7,  8'd2,  -8'd37,  8'd3,  
-8'd14,  8'd7,  -8'd15,  8'd18,  8'd50,  -8'd18,  8'd18,  
8'd18,  8'd24,  -8'd4,  8'd31,  -8'd3,  8'd3,  8'd9,  
-8'd1,  -8'd25,  -8'd34,  -8'd28,  8'd18,  -8'd2,  8'd0,  
-8'd7,  8'd3,  -8'd39,  -8'd17,  8'd15,  8'd10,  -8'd74,  
8'd7,  -8'd18,  -8'd6,  -8'd46,  8'd0,  -8'd48,  -8'd4,  
-8'd53,  8'd22,  -8'd38,  8'd25,  -8'd66,  -8'd17,  -8'd36,  
-8'd6,  -8'd41,  -8'd17,  -8'd45,  8'd9,  -8'd21,  8'd3,  

8'd27,  8'd51,  8'd52,  8'd27,  -8'd8,  8'd22,  -8'd21,  
-8'd12,  -8'd6,  -8'd8,  -8'd20,  8'd35,  8'd44,  8'd10,  
-8'd10,  8'd20,  8'd15,  8'd12,  -8'd15,  8'd34,  8'd7,  
8'd11,  -8'd22,  8'd41,  -8'd1,  8'd25,  -8'd7,  -8'd22,  
8'd24,  8'd51,  8'd4,  8'd5,  -8'd27,  8'd10,  -8'd17,  
8'd7,  -8'd21,  -8'd20,  -8'd24,  -8'd6,  -8'd14,  -8'd21,  
-8'd18,  8'd9,  8'd44,  -8'd33,  8'd0,  -8'd58,  8'd31,  
-8'd5,  -8'd19,  -8'd58,  -8'd5,  8'd17,  -8'd17,  -8'd30,  
-8'd5,  8'd45,  8'd0,  -8'd4,  -8'd27,  8'd13,  8'd7,  
8'd0,  -8'd24,  -8'd22,  -8'd26,  -8'd1,  8'd31,  8'd0,  
8'd34,  8'd16,  -8'd2,  -8'd15,  8'd40,  -8'd73,  8'd9,  
-8'd39,  -8'd10,  -8'd37,  -8'd58,  8'd32,  -8'd7,  -8'd17,  
8'd1,  8'd12,  -8'd10,  -8'd13,  8'd4,  8'd11,  -8'd11,  
-8'd40,  -8'd20,  -8'd2,  8'd7,  -8'd31,  8'd15,  -8'd39,  
-8'd30,  -8'd5,  8'd12,  -8'd101,  8'd59,  -8'd55,  -8'd22,  
8'd1,  -8'd17,  -8'd25,  8'd4,  8'd56,  8'd4,  -8'd6,  
-8'd15,  8'd34,  -8'd50,  -8'd37,  -8'd13,  8'd12,  -8'd19,  
-8'd6,  -8'd1,  8'd38,  -8'd9,  -8'd37,  8'd30,  -8'd71,  
8'd24,  -8'd17,  -8'd37,  8'd5,  8'd30,  -8'd6,  8'd19,  
8'd48,  -8'd10,  -8'd31,  8'd5,  8'd31,  -8'd10,  8'd4,  
8'd0,  8'd62,  8'd16,  8'd32,  8'd13,  8'd40,  8'd3,  
-8'd16,  8'd13,  8'd25,  -8'd4,  -8'd43,  -8'd29,  -8'd23,  
-8'd5,  8'd19,  -8'd21,  -8'd18,  8'd31,  8'd2,  8'd3,  
8'd41,  8'd11,  8'd50,  -8'd16,  8'd40,  -8'd7,  -8'd17,  
8'd24,  8'd49,  -8'd56,  -8'd25,  8'd23,  8'd24,  -8'd56,  
8'd14,  8'd27,  8'd37,  -8'd13,  8'd14,  8'd5,  8'd18,  
-8'd54,  8'd9,  8'd26,  8'd33,  -8'd31,  8'd42,  -8'd26,  
8'd55,  8'd8,  8'd8,  8'd5,  8'd61,  -8'd33,  -8'd59,  

-8'd9,  8'd4,  -8'd25,  -8'd35,  -8'd6,  -8'd12,  8'd7,  
-8'd20,  8'd7,  8'd19,  -8'd6,  -8'd10,  -8'd31,  -8'd2,  
8'd10,  8'd4,  -8'd2,  -8'd3,  8'd5,  -8'd18,  -8'd18,  
8'd11,  -8'd3,  -8'd50,  8'd0,  -8'd13,  8'd5,  8'd2,  
8'd12,  8'd13,  -8'd12,  8'd11,  -8'd11,  8'd19,  8'd6,  
-8'd7,  8'd0,  8'd12,  8'd30,  8'd16,  -8'd6,  -8'd5,  
8'd0,  8'd10,  -8'd42,  -8'd31,  8'd12,  8'd17,  -8'd25,  
-8'd29,  -8'd14,  8'd13,  -8'd15,  -8'd13,  -8'd21,  -8'd46,  
8'd24,  -8'd5,  8'd14,  -8'd20,  -8'd17,  8'd33,  8'd18,  
-8'd14,  -8'd36,  8'd52,  -8'd25,  -8'd10,  -8'd32,  8'd0,  
-8'd26,  -8'd3,  -8'd13,  -8'd20,  -8'd17,  8'd31,  8'd12,  
-8'd47,  8'd0,  -8'd17,  -8'd2,  -8'd11,  -8'd19,  -8'd44,  
-8'd6,  8'd15,  -8'd21,  -8'd14,  -8'd1,  8'd68,  -8'd13,  
-8'd79,  -8'd18,  8'd52,  -8'd21,  -8'd64,  -8'd16,  8'd37,  
-8'd5,  -8'd20,  8'd24,  8'd1,  -8'd6,  -8'd48,  8'd16,  
-8'd19,  8'd0,  -8'd27,  8'd38,  8'd41,  8'd3,  8'd14,  
8'd13,  8'd15,  8'd0,  8'd6,  8'd15,  -8'd9,  8'd12,  
-8'd10,  8'd55,  -8'd12,  8'd10,  -8'd32,  8'd33,  -8'd19,  
8'd28,  -8'd6,  8'd8,  8'd19,  8'd4,  -8'd4,  8'd1,  
8'd30,  8'd30,  -8'd13,  -8'd9,  8'd62,  -8'd10,  8'd32,  
8'd6,  -8'd6,  8'd7,  8'd16,  8'd8,  8'd0,  8'd6,  
-8'd1,  8'd31,  -8'd20,  8'd22,  8'd0,  -8'd21,  8'd16,  
-8'd3,  8'd17,  -8'd29,  8'd33,  8'd10,  8'd56,  -8'd36,  
8'd78,  8'd2,  8'd59,  8'd7,  8'd37,  -8'd39,  8'd5,  
8'd8,  -8'd3,  -8'd57,  -8'd45,  8'd15,  -8'd9,  -8'd78,  
8'd4,  -8'd18,  -8'd8,  -8'd24,  8'd0,  -8'd41,  -8'd19,  
-8'd17,  -8'd11,  -8'd41,  -8'd15,  8'd21,  8'd3,  -8'd45,  
-8'd16,  -8'd33,  8'd1,  8'd4,  8'd2,  -8'd8,  -8'd15,  

-8'd1,  -8'd19,  -8'd3,  8'd9,  8'd24,  -8'd16,  8'd15,  
-8'd12,  -8'd3,  -8'd19,  -8'd13,  -8'd11,  -8'd6,  -8'd14,  
8'd18,  -8'd6,  -8'd19,  -8'd2,  8'd12,  -8'd46,  -8'd6,  
-8'd27,  8'd23,  -8'd93,  8'd5,  -8'd30,  -8'd17,  -8'd25,  
-8'd25,  8'd0,  8'd22,  8'd0,  -8'd13,  8'd31,  8'd47,  
-8'd4,  -8'd22,  8'd27,  8'd40,  8'd32,  -8'd28,  8'd2,  
8'd28,  8'd23,  -8'd31,  -8'd28,  8'd16,  8'd8,  -8'd4,  
-8'd37,  8'd9,  -8'd8,  -8'd27,  -8'd39,  -8'd6,  -8'd46,  
8'd20,  -8'd31,  -8'd8,  8'd3,  8'd8,  8'd37,  8'd7,  
-8'd31,  -8'd37,  8'd55,  -8'd18,  -8'd51,  8'd10,  8'd50,  
8'd5,  -8'd18,  8'd40,  -8'd1,  8'd15,  -8'd15,  8'd19,  
-8'd30,  -8'd11,  -8'd24,  -8'd23,  -8'd38,  -8'd18,  -8'd14,  
8'd3,  8'd1,  -8'd22,  8'd12,  -8'd32,  8'd24,  -8'd46,  
-8'd56,  -8'd14,  8'd34,  -8'd16,  -8'd24,  8'd13,  8'd11,  
8'd9,  8'd5,  -8'd8,  8'd18,  -8'd4,  8'd14,  -8'd23,  
8'd8,  8'd1,  8'd10,  -8'd17,  -8'd31,  -8'd16,  -8'd3,  
8'd3,  8'd14,  8'd13,  8'd30,  -8'd25,  8'd38,  8'd1,  
8'd20,  -8'd58,  8'd21,  8'd1,  -8'd5,  -8'd50,  8'd30,  
-8'd2,  8'd38,  -8'd7,  8'd28,  -8'd6,  8'd26,  -8'd6,  
-8'd52,  8'd4,  -8'd1,  8'd12,  -8'd47,  8'd8,  -8'd9,  
-8'd10,  -8'd15,  -8'd9,  8'd0,  -8'd22,  8'd50,  8'd31,  
8'd1,  -8'd38,  8'd28,  8'd29,  -8'd9,  -8'd18,  8'd19,  
8'd19,  -8'd14,  8'd24,  -8'd10,  8'd9,  -8'd5,  8'd33,  
-8'd49,  8'd7,  -8'd11,  -8'd27,  -8'd66,  8'd0,  -8'd14,  
-8'd21,  -8'd48,  8'd54,  8'd71,  -8'd13,  8'd2,  8'd56,  
-8'd5,  8'd15,  8'd57,  8'd46,  -8'd4,  8'd0,  8'd52,  
8'd27,  -8'd28,  8'd15,  -8'd29,  -8'd24,  -8'd8,  8'd15,  
-8'd29,  8'd19,  -8'd16,  -8'd20,  -8'd37,  -8'd25,  -8'd14,  

8'd14,  8'd23,  8'd3,  8'd9,  -8'd6,  8'd11,  -8'd29,  
8'd0,  -8'd37,  -8'd17,  -8'd25,  -8'd10,  8'd4,  8'd0,  
-8'd29,  8'd6,  8'd8,  -8'd8,  -8'd32,  8'd0,  -8'd27,  
8'd2,  -8'd21,  8'd11,  8'd2,  8'd16,  -8'd31,  -8'd45,  
-8'd26,  8'd0,  8'd17,  8'd21,  8'd20,  -8'd5,  -8'd12,  
8'd22,  8'd14,  -8'd27,  -8'd36,  8'd43,  8'd30,  -8'd79,  
-8'd49,  -8'd4,  8'd53,  -8'd52,  -8'd30,  -8'd15,  8'd50,  
-8'd4,  -8'd2,  -8'd36,  8'd42,  8'd6,  8'd25,  8'd7,  
-8'd13,  -8'd4,  8'd3,  -8'd28,  -8'd10,  -8'd6,  -8'd8,  
8'd13,  8'd40,  -8'd33,  8'd8,  8'd26,  8'd25,  -8'd49,  
-8'd25,  -8'd52,  8'd57,  -8'd44,  8'd15,  -8'd38,  8'd30,  
-8'd17,  -8'd16,  -8'd72,  -8'd15,  -8'd8,  -8'd33,  -8'd27,  
-8'd19,  8'd3,  8'd29,  -8'd9,  8'd26,  8'd9,  8'd24,  
8'd20,  8'd50,  -8'd37,  8'd34,  8'd22,  -8'd12,  8'd17,  
8'd21,  8'd18,  8'd44,  -8'd19,  8'd29,  8'd0,  8'd24,  
8'd20,  8'd14,  -8'd7,  -8'd28,  8'd2,  8'd8,  -8'd4,  
8'd32,  -8'd13,  8'd0,  -8'd24,  8'd22,  -8'd9,  -8'd7,  
8'd3,  8'd7,  8'd19,  -8'd7,  -8'd15,  8'd1,  8'd10,  
-8'd15,  8'd29,  8'd1,  -8'd19,  8'd5,  8'd8,  -8'd8,  
-8'd15,  8'd0,  8'd22,  -8'd36,  8'd28,  -8'd26,  8'd2,  
-8'd49,  8'd0,  -8'd22,  -8'd22,  8'd4,  8'd26,  -8'd11,  
-8'd40,  -8'd9,  8'd12,  -8'd18,  -8'd59,  8'd0,  -8'd93,  
-8'd43,  -8'd17,  -8'd14,  -8'd85,  8'd6,  8'd3,  -8'd7,  
8'd2,  8'd15,  -8'd3,  -8'd19,  8'd29,  8'd5,  -8'd2,  
-8'd46,  8'd17,  -8'd2,  -8'd25,  -8'd4,  -8'd7,  8'd18,  
-8'd22,  8'd24,  -8'd75,  8'd13,  8'd11,  8'd3,  -8'd55,  
8'd3,  8'd13,  8'd15,  8'd15,  -8'd8,  8'd30,  8'd20,  
-8'd1,  -8'd29,  8'd26,  -8'd9,  8'd30,  8'd13,  -8'd8,  

8'd19,  8'd20,  -8'd15,  -8'd18,  -8'd41,  8'd9,  -8'd33,  
-8'd12,  -8'd6,  8'd1,  8'd0,  -8'd25,  -8'd18,  -8'd3,  
8'd3,  -8'd21,  8'd8,  8'd11,  8'd13,  8'd23,  8'd2,  
-8'd12,  8'd10,  8'd24,  8'd6,  8'd9,  -8'd10,  8'd25,  
-8'd18,  -8'd10,  -8'd34,  -8'd21,  -8'd13,  -8'd2,  -8'd19,  
-8'd15,  8'd0,  -8'd7,  -8'd11,  8'd1,  -8'd11,  -8'd1,  
8'd7,  -8'd36,  -8'd8,  8'd35,  8'd8,  -8'd2,  8'd5,  
8'd46,  8'd41,  -8'd2,  8'd18,  8'd24,  8'd15,  -8'd6,  
-8'd61,  8'd4,  8'd7,  -8'd42,  -8'd2,  -8'd62,  -8'd35,  
8'd15,  8'd3,  -8'd42,  8'd23,  8'd17,  -8'd10,  8'd26,  
8'd10,  -8'd32,  -8'd101,  8'd42,  -8'd14,  8'd2,  -8'd93,  
8'd81,  -8'd6,  8'd15,  8'd14,  8'd52,  -8'd20,  8'd57,  
-8'd2,  -8'd6,  -8'd15,  -8'd6,  8'd1,  -8'd39,  8'd19,  
8'd11,  -8'd13,  8'd0,  8'd15,  8'd31,  -8'd36,  8'd13,  
8'd3,  8'd5,  -8'd76,  8'd2,  -8'd17,  8'd25,  -8'd72,  
8'd33,  -8'd35,  8'd0,  -8'd26,  8'd59,  -8'd58,  -8'd15,  
-8'd3,  8'd33,  -8'd1,  8'd3,  -8'd50,  8'd57,  -8'd14,  
8'd21,  -8'd56,  8'd43,  -8'd10,  8'd17,  -8'd20,  8'd10,  
8'd4,  8'd10,  -8'd1,  8'd9,  8'd8,  8'd11,  8'd1,  
-8'd59,  8'd3,  8'd8,  8'd13,  -8'd11,  8'd18,  -8'd22,  
-8'd14,  -8'd3,  -8'd9,  -8'd20,  -8'd22,  8'd50,  8'd4,  
8'd9,  -8'd31,  8'd29,  8'd19,  8'd11,  8'd10,  8'd20,  
8'd16,  -8'd24,  8'd24,  8'd14,  8'd9,  -8'd7,  8'd36,  
-8'd32,  8'd17,  8'd0,  8'd35,  -8'd19,  8'd26,  8'd9,  
-8'd16,  -8'd2,  8'd2,  -8'd39,  -8'd30,  -8'd3,  8'd15,  
-8'd31,  -8'd2,  8'd23,  8'd33,  -8'd22,  -8'd8,  8'd59,  
8'd27,  -8'd13,  8'd16,  8'd22,  8'd3,  -8'd5,  8'd35,  
8'd29,  -8'd16,  -8'd27,  8'd27,  8'd27,  8'd33,  8'd34,  

-8'd22,  8'd1,  8'd30,  8'd37,  8'd13,  -8'd6,  8'd31,  
8'd38,  8'd52,  -8'd10,  8'd25,  8'd26,  8'd17,  8'd0,  
-8'd19,  8'd22,  8'd29,  8'd8,  8'd20,  8'd5,  8'd7,  
8'd24,  8'd37,  8'd34,  8'd10,  -8'd1,  8'd33,  8'd14,  
8'd1,  -8'd2,  -8'd9,  -8'd31,  8'd8,  -8'd14,  8'd10,  
8'd8,  -8'd5,  -8'd41,  -8'd34,  -8'd38,  8'd45,  -8'd6,  
-8'd32,  -8'd57,  8'd0,  8'd2,  -8'd24,  -8'd34,  -8'd14,  
8'd22,  -8'd6,  8'd22,  8'd6,  -8'd22,  -8'd1,  8'd43,  
-8'd18,  -8'd21,  -8'd8,  -8'd24,  8'd21,  -8'd31,  -8'd16,  
-8'd15,  8'd33,  -8'd18,  8'd6,  -8'd13,  8'd19,  -8'd17,  
-8'd18,  -8'd78,  -8'd21,  8'd48,  -8'd35,  -8'd40,  -8'd43,  
8'd51,  -8'd29,  8'd30,  -8'd30,  -8'd5,  -8'd4,  -8'd19,  
-8'd76,  -8'd33,  8'd3,  8'd2,  8'd18,  -8'd44,  -8'd6,  
8'd1,  8'd38,  -8'd63,  -8'd14,  -8'd36,  8'd13,  8'd12,  
8'd18,  -8'd38,  -8'd32,  8'd44,  8'd7,  8'd4,  -8'd11,  
8'd5,  8'd0,  8'd19,  8'd30,  -8'd53,  8'd18,  8'd24,  
-8'd21,  -8'd31,  -8'd26,  -8'd38,  -8'd9,  -8'd90,  -8'd6,  
8'd26,  8'd18,  -8'd55,  8'd13,  8'd45,  8'd4,  -8'd13,  
8'd30,  8'd16,  8'd3,  -8'd5,  8'd9,  8'd21,  8'd24,  
-8'd20,  8'd24,  -8'd4,  8'd16,  -8'd26,  8'd28,  8'd2,  
-8'd46,  -8'd16,  -8'd38,  -8'd33,  8'd11,  -8'd60,  -8'd13,  
8'd20,  -8'd21,  -8'd35,  8'd22,  8'd37,  -8'd24,  8'd11,  
8'd32,  8'd47,  8'd1,  8'd8,  8'd18,  8'd20,  -8'd1,  
8'd0,  -8'd20,  8'd9,  8'd27,  -8'd2,  -8'd16,  -8'd7,  
-8'd67,  -8'd9,  -8'd9,  -8'd27,  -8'd40,  -8'd3,  -8'd25,  
-8'd70,  -8'd5,  -8'd1,  -8'd54,  -8'd31,  -8'd46,  8'd5,  
-8'd48,  -8'd33,  -8'd44,  -8'd9,  -8'd31,  -8'd25,  -8'd48,  
-8'd9,  -8'd4,  -8'd1,  -8'd45,  -8'd4,  -8'd47,  -8'd23,  

-8'd14,  8'd24,  -8'd11,  -8'd15,  8'd12,  8'd35,  8'd24,  
8'd32,  -8'd28,  8'd7,  -8'd25,  8'd6,  -8'd11,  8'd17,  
-8'd17,  -8'd35,  -8'd12,  8'd1,  -8'd11,  -8'd72,  -8'd30,  
-8'd4,  -8'd59,  -8'd39,  -8'd66,  8'd18,  -8'd47,  -8'd4,  
8'd50,  8'd9,  8'd5,  -8'd19,  8'd12,  8'd17,  8'd3,  
8'd19,  8'd0,  8'd42,  8'd23,  8'd36,  -8'd35,  -8'd2,  
8'd4,  8'd8,  8'd6,  8'd20,  -8'd10,  -8'd11,  8'd16,  
8'd2,  -8'd11,  -8'd29,  -8'd4,  -8'd2,  -8'd17,  -8'd58,  
8'd6,  8'd25,  8'd8,  8'd24,  -8'd17,  8'd32,  8'd41,  
8'd28,  -8'd24,  8'd9,  8'd31,  8'd10,  -8'd14,  8'd24,  
8'd8,  8'd31,  8'd29,  8'd0,  8'd37,  8'd42,  8'd21,  
-8'd14,  8'd13,  -8'd32,  -8'd22,  -8'd13,  8'd13,  -8'd46,  
8'd15,  8'd19,  8'd16,  8'd14,  -8'd1,  8'd27,  8'd20,  
-8'd24,  8'd27,  8'd9,  -8'd48,  -8'd73,  8'd3,  -8'd4,  
-8'd61,  -8'd51,  8'd12,  -8'd17,  -8'd1,  -8'd26,  8'd23,  
8'd54,  8'd3,  -8'd2,  -8'd11,  8'd6,  -8'd22,  -8'd48,  
-8'd25,  8'd17,  -8'd26,  -8'd22,  8'd14,  8'd3,  -8'd24,  
-8'd33,  -8'd8,  -8'd4,  -8'd1,  -8'd15,  8'd15,  -8'd9,  
-8'd36,  -8'd38,  8'd12,  -8'd16,  8'd25,  -8'd15,  -8'd10,  
-8'd4,  8'd5,  8'd39,  -8'd59,  8'd19,  -8'd32,  -8'd20,  
8'd6,  8'd36,  -8'd12,  -8'd12,  8'd11,  8'd6,  8'd4,  
-8'd43,  8'd16,  -8'd21,  -8'd38,  -8'd54,  8'd10,  -8'd83,  
-8'd31,  -8'd9,  -8'd20,  -8'd62,  -8'd19,  -8'd31,  -8'd37,  
-8'd33,  -8'd26,  -8'd31,  -8'd60,  8'd4,  -8'd82,  -8'd52,  
8'd24,  8'd33,  8'd42,  8'd3,  8'd46,  -8'd3,  8'd20,  
8'd22,  8'd16,  8'd6,  8'd19,  8'd35,  8'd17,  8'd7,  
8'd15,  8'd24,  8'd32,  -8'd10,  8'd38,  8'd4,  -8'd23,  
8'd38,  8'd15,  -8'd7,  -8'd4,  8'd13,  -8'd19,  -8'd41,  

-8'd40,  -8'd50,  -8'd63,  -8'd37,  -8'd4,  -8'd20,  8'd10,  
8'd0,  8'd8,  8'd29,  -8'd11,  -8'd17,  -8'd9,  8'd0,  
-8'd6,  8'd2,  8'd19,  8'd10,  8'd0,  8'd13,  -8'd9,  
-8'd8,  -8'd3,  -8'd20,  8'd4,  -8'd26,  8'd14,  8'd18,  
-8'd26,  -8'd31,  -8'd22,  -8'd3,  8'd3,  -8'd21,  -8'd18,  
-8'd6,  8'd0,  8'd3,  -8'd8,  -8'd14,  8'd21,  8'd23,  
-8'd7,  -8'd13,  -8'd10,  8'd3,  -8'd20,  8'd40,  -8'd12,  
8'd16,  -8'd4,  8'd19,  -8'd15,  -8'd8,  8'd7,  8'd37,  
-8'd8,  -8'd28,  -8'd2,  8'd34,  8'd13,  -8'd9,  8'd2,  
8'd31,  -8'd14,  -8'd10,  -8'd16,  8'd53,  -8'd29,  -8'd2,  
-8'd10,  8'd33,  8'd3,  -8'd3,  8'd0,  -8'd3,  8'd30,  
8'd7,  8'd11,  8'd13,  8'd36,  -8'd20,  8'd10,  -8'd18,  
-8'd14,  -8'd50,  -8'd5,  8'd0,  8'd5,  -8'd28,  8'd10,  
8'd6,  -8'd20,  -8'd15,  -8'd20,  8'd48,  8'd21,  -8'd16,  
8'd23,  8'd42,  8'd5,  8'd6,  8'd0,  -8'd22,  -8'd9,  
8'd26,  -8'd26,  8'd27,  8'd1,  -8'd58,  -8'd14,  8'd45,  
-8'd41,  -8'd36,  -8'd3,  -8'd5,  8'd10,  8'd3,  8'd8,  
-8'd30,  8'd51,  -8'd16,  -8'd16,  -8'd18,  -8'd13,  -8'd27,  
-8'd18,  8'd26,  -8'd32,  8'd14,  -8'd46,  8'd25,  -8'd26,  
-8'd9,  -8'd12,  8'd20,  8'd9,  -8'd42,  -8'd12,  -8'd17,  
-8'd15,  -8'd33,  8'd2,  -8'd21,  8'd25,  -8'd51,  -8'd4,  
8'd2,  -8'd7,  -8'd35,  8'd15,  8'd11,  -8'd5,  -8'd3,  
8'd28,  8'd12,  8'd19,  8'd19,  8'd8,  8'd4,  8'd27,  
-8'd38,  8'd2,  -8'd8,  -8'd21,  -8'd46,  8'd25,  8'd15,  
8'd6,  -8'd68,  -8'd67,  -8'd83,  8'd5,  -8'd63,  -8'd34,  
8'd3,  -8'd25,  -8'd86,  -8'd7,  8'd9,  -8'd3,  -8'd50,  
8'd4,  8'd2,  -8'd19,  -8'd49,  -8'd20,  -8'd5,  8'd18,  
-8'd56,  -8'd34,  -8'd2,  -8'd42,  -8'd31,  -8'd12,  8'd0,  

-8'd14,  -8'd30,  -8'd28,  -8'd34,  -8'd53,  -8'd25,  8'd1,  
-8'd28,  -8'd13,  8'd7,  8'd18,  -8'd18,  8'd4,  -8'd2,  
-8'd1,  -8'd74,  -8'd22,  -8'd30,  -8'd7,  -8'd42,  8'd4,  
-8'd19,  8'd1,  -8'd93,  -8'd36,  -8'd52,  -8'd57,  -8'd6,  
-8'd74,  -8'd41,  -8'd20,  -8'd25,  8'd6,  8'd0,  -8'd1,  
-8'd48,  -8'd15,  8'd27,  -8'd6,  -8'd65,  8'd1,  8'd60,  
8'd26,  8'd12,  -8'd28,  8'd18,  8'd26,  8'd7,  -8'd46,  
-8'd8,  -8'd5,  8'd21,  -8'd52,  -8'd25,  -8'd20,  -8'd47,  
-8'd13,  8'd0,  -8'd3,  8'd2,  8'd7,  -8'd5,  -8'd4,  
8'd2,  8'd48,  8'd0,  -8'd34,  -8'd2,  8'd1,  8'd5,  
-8'd16,  8'd4,  8'd4,  8'd29,  -8'd4,  8'd14,  -8'd6,  
-8'd22,  -8'd6,  8'd11,  -8'd30,  -8'd37,  -8'd1,  -8'd26,  
8'd8,  -8'd50,  -8'd6,  8'd31,  8'd6,  -8'd54,  8'd0,  
8'd27,  -8'd14,  -8'd26,  8'd36,  8'd43,  8'd7,  8'd29,  
8'd50,  8'd11,  8'd16,  -8'd18,  8'd15,  8'd18,  8'd16,  
-8'd73,  8'd20,  -8'd11,  -8'd39,  -8'd61,  8'd11,  -8'd26,  
8'd9,  -8'd54,  -8'd10,  8'd2,  -8'd9,  -8'd44,  8'd10,  
8'd34,  -8'd55,  8'd42,  8'd13,  8'd32,  -8'd13,  8'd33,  
-8'd54,  -8'd12,  8'd9,  -8'd36,  -8'd30,  -8'd18,  8'd1,  
-8'd102,  -8'd12,  -8'd31,  -8'd45,  -8'd24,  8'd2,  -8'd31,  
-8'd18,  -8'd43,  8'd1,  -8'd7,  8'd7,  8'd16,  8'd3,  
-8'd19,  -8'd12,  8'd32,  -8'd41,  -8'd28,  8'd6,  -8'd1,  
-8'd54,  -8'd31,  -8'd10,  -8'd24,  -8'd2,  -8'd17,  8'd17,  
-8'd21,  -8'd5,  -8'd3,  8'd18,  8'd13,  8'd15,  -8'd8,  
-8'd3,  8'd7,  8'd38,  8'd27,  8'd28,  8'd16,  8'd4,  
-8'd14,  8'd31,  8'd19,  8'd1,  -8'd10,  8'd6,  -8'd44,  
8'd16,  -8'd2,  8'd6,  -8'd40,  8'd16,  8'd26,  8'd38,  
-8'd22,  8'd13,  8'd7,  -8'd15,  -8'd17,  8'd3,  8'd10



};
	always @(posedge clk or negedge rst_n)
		if (!rst_n)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule



